package tb_os_specific_only;
    parameter string myLeds = "/Volumes/RAM_Disk_4G/tmpFifo/myLeds";
    parameter string mySegDispllay = "/Volumes/RAM_Disk_4G/tmpFifo/my7SegDispllay";
    parameter string mySw = "/Volumes/RAM_Disk_4G/tmpFifo/mySw";
    parameter string myBtns = "/Volumes/RAM_Disk_4G/tmpFifo/myBtns";
endpackage