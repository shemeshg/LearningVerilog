`timescale 1ns / 10ps
module select_btn_action (
    input  word_t SW,
    output word_t LED,
    input  wire   rst,
    input  wire   clk,
    input  wire   BTNC,
    input  wire   BTNU,
    input  wire   BTNL,
    input  wire   BTNR,
    input  wire   BTND,
    output int    calc_displayed,
    output logic  isEdit
);
  import types_pkg::*;

  // *** IMPORTANT FIX ***
  // total must be SIGNED or subtraction will wrap around
  logic signed [BITS-1:0] total;

  // LED mirrors switches
  always_comb begin
    LED = SW;
    calc_displayed = isEdit ? int'(SW) : int'(total);
  end

  // Edge detectors
  logic rise_u, rise_d, rise_r, rise_l, rise_c;

  edge_detect ed_u (.clk(clk), .rst(rst), .sig(BTNU), .rise(rise_u));
  edge_detect ed_d (.clk(clk), .rst(rst), .sig(BTND), .rise(rise_d));
  edge_detect ed_r (.clk(clk), .rst(rst), .sig(BTNR), .rise(rise_r));
  edge_detect ed_l (.clk(clk), .rst(rst), .sig(BTNL), .rise(rise_l));
  edge_detect ed_c (.clk(clk), .rst(rst), .sig(BTNC), .rise(rise_c));

  // Divider
  logic        div_start, div_done;
  logic        div_busy;
  logic [BITS-1:0] div_quotient, div_remainder;

  divider_nr u_divider (
      .clk(clk),
      .reset(rst),
      .start(div_start),
      .dividend(total),
      .divisor(SW),
      .done(div_done),
      .quotient(div_quotient),
      .remainder(div_remainder)
  );

  // Main state logic
  always_ff @(posedge clk) begin
    if (rst) begin
      total     <= '0;
      isEdit    <= 1;
      div_start <= 0;
      div_busy  <= 0;
    end else begin
      // defaults
      div_start <= 0;

      // arithmetic operations
      if (rise_u) total <= total + $signed(SW);
      if (rise_d) total <= total - $signed(SW);
      if (rise_r) total <= total * $signed(SW);

      // toggle edit mode
      if (rise_c) isEdit <= ~isEdit;

      // start division
      if (rise_l && !div_busy && SW != 0) begin
        div_start <= 1;
        div_busy  <= 1;
      end

      // division result
      if (div_done) begin
        total    <= $signed(div_quotient);
        div_busy <= 0;
      end
    end
  end

endmodule
