import types_pkg::*;

module seg_display (
    input display_t display,
    input wire CLK100MHZ,
    input wire CPU_RESET,
    input word_t SW,
    output word_t  LED,
    input wire                     BTNC,
    input wire                     BTNU,
    input wire                     BTNL,
    input wire                     BTNR,
    input wire                     BTND,      
    output word_t AN,
    output wire   CA,
    output wire   CB,
    output wire   CC,
    output wire   CD,
    output wire   CE,
    output wire   CF,
    output wire   CG,
    output wire   DP
);



endmodule
