package tb_os_specific_only;
    parameter string myLeds = "/dev/shm/myLeds";
    parameter string mySegDispllay = "/dev/shm/my7SegDispllay";
    parameter string mySw = "/dev/shm/mySw";
    parameter string myBtns = "/dev/shm/myBtns";
endpackage