import types_pkg::*;

module seg_display (
    input display_t display,
    input wire CPU_RESET,
    input wire CLOCK,
    output word_t AN,
    output wire   CA,
    output wire   CB,
    output wire   CC,
    output wire   CD,
    output wire   CE,
    output wire   CF,
    output wire   CG,
    output wire   DP
);



endmodule
